class transaction;
 
  randc reg[7:0] A,B;
  reg[3:0] ALU_Sel;
  reg clk;
  logic [7:0] ALU_Out;
  logic CarryOut;
           
endclass
